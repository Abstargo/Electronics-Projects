CircuitMaker Text
5.6
Probes: 1
Vs
Transient Analysis
0 246 95 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1022 385
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
51 C:\LOGICIEL DE SIMULATION\CIRCUITMAKER 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1190 489
9961490 0
0
6 Title:
5 Name:
0
0
0
14
2 +V
167 225 43 0 1 3
0 5
0
0 0 54112 0
3 10V
-11 -22 10 -14
3 Vss
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6316 0 0
2
5.90027e-315 0
0
2 +V
167 222 164 0 1 3
0 4
0
0 0 54112 180
4 -10V
3 -2 31 6
3 Vdd
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8734 0 0
2
5.90027e-315 5.26354e-315
0
5 SAVE-
218 96 160 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 C
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
7988 0 0
2
5.90027e-315 5.30499e-315
0
5 SAVE-
218 106 85 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3217 0 0
2
5.90027e-315 5.32571e-315
0
5 SAVE-
218 225 94 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3965 0 0
2
5.90027e-315 5.34643e-315
0
9 Terminal~
194 247 84 0 1 3
0 2
0
0 0 49504 0
2 Vs
-6 -13 8 -5
2 T1
-7 -32 7 -24
0
3 Vs;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8239 0 0
2
5.90027e-315 5.3568e-315
0
11 Signal Gen~
195 46 165 0 64 64
0 6 3 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1120403456 0 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 100 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -500m/500mV
-39 -30 38 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 500m 100 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
828 0 0
2
5.90027e-315 5.36716e-315
0
8 Battery~
219 148 164 0 2 5
0 7 3
0
0 0 864 0
5 0.75V
6 -2 41 6
2 V0
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6187 0 0
2
5.90027e-315 5.37752e-315
0
7 Ground~
168 93 187 0 1 3
0 3
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7107 0 0
2
5.90027e-315 5.38788e-315
0
7 Ground~
168 280 141 0 1 3
0 3
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6433 0 0
2
5.90027e-315 5.39306e-315
0
7 Ground~
168 94 122 0 1 3
0 3
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8559 0 0
2
5.90027e-315 5.39824e-315
0
11 Signal Gen~
195 47 89 0 19 64
0 8 3 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1084227584
20
1 10000 0 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 -5/5V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 5 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3674 0 0
2
5.90027e-315 5.40342e-315
0
7 Ground~
168 148 224 0 1 3
0 3
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5697 0 0
2
5.90027e-315 5.4086e-315
0
6 AD633~
219 185 103 0 8 17
0 8 3 6 7 4 3 2 5
0
0 0 4928 0
5 AD633
-17 -37 18 -29
2 U1
-6 -47 8 -39
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 14346004
88 0 0 256 1 1 0 0
1 U
3805 0 0
2
5.90027e-315 5.41378e-315
0
11
5 1 4 0 0 8320 0 14 2 0 0 3
218 112
222 112
222 149
8 1 5 0 0 4224 0 14 1 0 0 3
218 85
218 52
225 52
6 1 3 0 0 4224 0 14 10 0 0 3
218 103
280 103
280 135
1 7 2 0 0 8320 0 6 14 0 0 3
247 93
247 94
218 94
2 1 3 0 0 0 0 7 9 0 0 3
77 170
93 170
93 181
3 1 6 0 0 8320 0 14 7 0 0 4
152 103
117 103
117 160
77 160
2 1 3 0 0 0 0 8 13 0 0 2
148 175
148 218
4 1 7 0 0 8320 0 14 8 0 0 3
152 112
148 112
148 151
2 0 3 0 0 0 0 14 0 0 10 2
152 94
94 94
2 1 3 0 0 0 0 12 11 0 0 3
78 94
94 94
94 116
1 1 8 0 0 4224 0 14 12 0 0 4
152 85
86 85
86 84
78 84
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.05 0.0001 0.0001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
