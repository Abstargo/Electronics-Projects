CircuitMaker Text
5.6
Probes: 13
V2_1
AC Analysis
2 124 225 16776960
V2_1
DC Sweep
2 124 225 16776960
V2_1
Operating Point
2 124 225 16776960
V2_1
Transient Analysis
2 124 225 16776960
V1_1
AC Analysis
1 130 130 65535
V1_1
DC Sweep
1 130 130 65535
V1_1
Operating Point
1 130 130 65535
V1_1
Transient Analysis
1 130 130 65535
Vs
AC Analysis
0 242 169 65280
Vs
DC Sweep
0 242 169 65280
Vs
Operating Point
0 242 169 65280
Vs
Transient Analysis
0 242 169 65280
Vs
Fourier Analysis
0 250 167 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1022 385
7 5.000 V
7 5.000 V
3 GND
30000 4
24 100 0 1 0
20 Package,Description,
51 C:\LOGICIEL DE SIMULATION\CIRCUITMAKER 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1190 489
9961490 0
0
6 Title:
5 Name:
0
0
0
9
9 Terminal~
194 268 157 0 1 3
0 2
0
0 0 49520 0
2 Vs
-7 -22 7 -14
2 T1
-7 -32 7 -24
0
3 Vs;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7804 0 0
2
5.89339e-315 0
0
11 Signal Gen~
195 61 136 0 64 64
0 4 3 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1189765120 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 30000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
30 %D %1 %2 DC 0 SIN(0 1 30k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5523 0 0
2
44663.7 0
0
5 SAVE-
218 124 225 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 C
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3330 0 0
2
44663.7 1
0
5 SAVE-
218 130 130 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3465 0 0
2
44663.7 2
0
5 SAVE-
218 242 169 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
8396 0 0
2
44663.7 3
0
7 Ground~
168 94 255 0 1 3
0 3
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3685 0 0
2
44663.7 4
0
11 Signal Gen~
195 61 230 0 64 64
0 5 3 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1189765120 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 30000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V2
-7 -40 7 -32
0
0
30 %D %1 %2 DC 0 SIN(0 1 30k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7849 0 0
2
44663.7 5
0
7 Ground~
168 100 172 0 1 3
0 3
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6343 0 0
2
5.89339e-315 0
0
11 multiplier~
219 188 169 0 3 7
0 4 5 2
0
0 0 50000 0
4 MULT
-7 -31 21 -23
2 U1
0 -41 14 -33
0
0
16 %D [%1 %2] %3 %M
0
15 type:multiplier
0
7

0 0 0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
7376 0 0
2
5.89339e-315 5.30499e-315
0
5
1 3 2 0 0 8320 0 1 9 0 0 3
268 166
268 169
226 169
2 1 3 0 0 8320 0 2 8 0 0 3
92 141
100 141
100 166
1 1 4 0 0 4224 0 2 9 0 0 4
92 131
156 131
156 160
164 160
1 2 5 0 0 4224 0 7 9 0 0 4
92 225
156 225
156 178
164 178
1 2 3 0 0 0 0 6 7 0 0 3
94 249
94 235
92 235
0
0
49 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.0001667 6.667e-07 2e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1212 2259520 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
0 0 0 0 0 0
12409 0
4 1 0.1
1
113 28
0 5 0 0 1	10 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
