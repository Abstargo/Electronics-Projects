CircuitMaker Text
5.6
Probes: 11
Vs
AC Analysis
0 237 169 65280
Vs
DC Sweep
0 237 169 65280
Vs
Fourier Analysis
0 237 169 65280
V2_1
AC Analysis
2 123 186 16776960
V2_1
DC Sweep
2 123 186 16776960
V2_1
Fourier Analysis
2 123 186 16776960
V1_1
AC Analysis
1 124 115 65535
V1_1
DC Sweep
1 124 115 65535
V1_1
Fourier Analysis
1 124 115 65535
Vs
Operating Point
0 241 169 65280
Vs
Transient Analysis
0 234 168 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1022 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
51 C:\LOGICIEL DE SIMULATION\CIRCUITMAKER 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1190 489
9961490 0
0
6 Title:
5 Name:
0
0
0
9
9 V Source~
197 58 213 0 2 5
0 4 3
0
0 0 17264 0
2 3V
16 0 30 8
2 V2
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
972 0 0
2
44663.7 0
0
5 SAVE-
218 237 169 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3472 0 0
2
44663.7 1
0
9 Terminal~
194 270 156 0 1 3
0 2
0
0 0 49520 0
2 Vs
-7 -22 7 -14
2 T1
-7 -32 7 -24
0
3 Vs;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9998 0 0
2
44663.7 2
0
9 V Source~
197 56 137 0 2 5
0 5 3
0
0 0 17264 0
2 0V
16 0 30 8
2 V1
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3536 0 0
2
44663.7 3
0
5 SAVE-
218 123 186 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 C
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
4597 0 0
2
44663.7 4
0
5 SAVE-
218 124 115 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3835 0 0
2
44663.7 5
0
7 Ground~
168 92 256 0 1 3
0 3
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
44663.7 6
0
7 Ground~
168 91 173 0 1 3
0 3
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
5.90027e-315 0
0
11 multiplier~
219 188 168 0 3 7
0 5 4 2
0
0 0 50000 0
4 MULT
-7 -31 21 -23
2 U1
0 -41 14 -33
0
0
16 %D [%1 %2] %3 %M
0
15 type:multiplier
0
7

0 0 0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
9323 0 0
2
5.90027e-315 5.26354e-315
0
5
2 1 3 0 0 8192 0 1 7 0 0 4
58 234
58 241
92 241
92 250
1 2 4 0 0 8320 0 1 9 0 0 5
58 192
58 186
156 186
156 177
164 177
3 1 2 0 0 4224 0 9 3 0 0 3
226 168
270 168
270 165
1 2 3 0 0 8320 0 8 4 0 0 4
91 167
91 164
56 164
56 158
1 1 5 0 0 8320 0 4 9 0 0 5
56 116
56 115
156 115
156 159
164 159
0
0
16 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.0001667 6.667e-07 6.667e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1212 2259520 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
0 0 0 0 0 0
12409 0
4 1 0.1
1
113 28
0 5 0 0 1	10 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
