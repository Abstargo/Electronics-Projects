CircuitMaker Text
5.6
Probes: 13
Vs
AC Analysis
0 277 125 65280
Vs
DC Sweep
0 277 125 65280
Vs
Operating Point
0 277 125 65280
Vs
Fourier Analysis
0 277 125 65280
V1_1
AC Analysis
2 158 182 16776960
V1_1
DC Sweep
2 158 182 16776960
V1_1
Operating Point
2 158 182 16776960
V1_1
Fourier Analysis
2 158 182 16776960
V2_1
AC Analysis
1 154 117 65535
V2_1
DC Sweep
1 154 117 65535
V2_1
Operating Point
1 154 117 65535
V2_1
Fourier Analysis
1 154 117 65535
Vs
Transient Analysis
0 301 118 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1022 385
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
51 C:\LOGICIEL DE SIMULATION\CIRCUITMAKER 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1190 489
9961490 0
0
6 Title:
5 Name:
0
0
0
15
10 Capacitor~
219 764 246 0 2 5
0 2 5
0
0 0 848 90
3 1�F
11 0 32 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5219 0 0
2
5.898e-315 0
0
6 Diode~
219 475 220 0 2 5
0 3 6
0
0 0 848 0
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3795 0 0
2
5.898e-315 0
0
10 Capacitor~
219 626 236 0 2 5
0 2 6
0
0 0 848 90
5 220nF
5 0 40 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3637 0 0
2
5.898e-315 0
0
7 Ground~
168 509 294 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3226 0 0
2
5.898e-315 0
0
5 SAVE-
218 277 125 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
6966 0 0
2
44663.7 0
0
5 SAVE-
218 158 182 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 C
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
9796 0 0
2
44663.7 1
0
5 SAVE-
218 154 117 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
5952 0 0
2
44663.7 2
0
9 Terminal~
194 301 107 0 1 3
0 3
0
0 0 49520 0
2 Vs
-7 -22 7 -14
2 T1
-7 -32 7 -24
0
3 Vs;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3649 0 0
2
44663.7 3
0
7 Ground~
168 98 210 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3716 0 0
2
5.898e-315 0
0
7 Ground~
168 103 137 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4797 0 0
2
5.898e-315 5.26354e-315
0
11 Signal Gen~
195 67 187 0 19 64
0 7 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1157070848 0 1067030938
20
0 1980 0 1.2 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -1.2/1.2V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
34 %D %1 %2 DC 0 SIN(0 1.2 1.98k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4681 0 0
2
5.898e-315 5.30499e-315
0
11 Signal Gen~
195 68 122 0 19 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1056964608 1157234688 0 1069547520
20
0.5 2000 0 1.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -1.5/1.5V
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
41 %D %1 %2 DC 0 SIN(0 1.5 2k 0 0) AC 500m 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9730 0 0
2
5.898e-315 5.32571e-315
0
7 summer~
219 223 126 0 3 7
0 8 7 3
0
0 0 50000 0
3 SUM
-4 -31 17 -23
2 U1
0 -41 14 -33
0
0
16 %D [%1 %2] %3 %M
0
11 type:summer
0
7

0 0 0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
9874 0 0
2
5.898e-315 5.34643e-315
0
9 Resistor~
219 708 214 0 2 5
0 6 5
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
364 0 0
2
5.898e-315 0
0
9 Resistor~
219 571 236 0 3 5
0 2 6 -1
0
0 0 880 90
3 10k
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3656 0 0
2
5.898e-315 0
0
14
0 0 4 0 0 4224 0 0 0 0 0 2
780 411
780 401
1 0 2 0 0 8320 0 1 0 0 7 3
764 255
764 260
626 260
2 2 5 0 0 4224 0 14 1 0 0 3
726 214
764 214
764 237
1 0 6 0 0 4096 0 14 0 0 8 2
690 214
626 214
1 1 3 0 0 4224 0 2 8 0 0 3
465 220
301 220
301 116
0 1 2 0 0 0 0 0 4 7 0 4
571 262
571 280
509 280
509 288
1 1 2 0 0 0 0 3 15 0 0 4
626 245
626 262
571 262
571 254
2 2 6 0 0 0 0 15 3 0 0 4
571 218
571 214
626 214
626 227
2 2 6 0 0 4224 0 2 15 0 0 5
485 220
563 220
563 210
571 210
571 218
1 3 3 0 0 0 0 8 13 0 0 3
301 116
301 126
261 126
1 2 7 0 0 4224 0 11 13 0 0 4
98 182
181 182
181 135
199 135
1 1 8 0 0 4224 0 12 13 0 0 2
99 117
199 117
1 2 2 0 0 0 0 9 11 0 0 2
98 204
98 192
1 2 2 0 0 0 0 10 12 0 0 3
103 131
103 127
99 127
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.15 0.0005 1.01e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1212 2259520 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
0 0 0 0 0 0
12409 0
4 1 0.1
1
113 28
0 5 0 0 1	16 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
